//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 (64-bit)
//Part Number: GW1NR-UV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Mon Sep  8 20:11:19 2025

module rom (dout, clk, oce, ce, reset, ad);

output wire [7:0] dout;
input wire clk;
input wire oce;
input wire ce;
input wire reset;
input wire [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hA9FF65018D0060A0FFA2FFCAD0FD88D0F84C0280B195817E0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000001038BCFFBC381000383A9FFF9F3A3800081C3E7F3E1C08;
defparam prom_inst_0.INIT_RAM_02 = 256'h0F077FFD8888F870000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h995A3CE7E73C5A993F7F6505057FFFC00000000000000000004E5FF1F15F4E00;
defparam prom_inst_0.INIT_RAM_04 = 256'h005F5F00005F5F00002466FFFF662400007F3E3E1C1C08080008081C1C3E3E7F;
defparam prom_inst_0.INIT_RAM_05 = 256'h8094B6FFFFB694800070707070707000020359FDA5A5BFDA7F7F017F7F090F06;
defparam prom_inst_0.INIT_RAM_06 = 256'h000808082A3E1C0800081C3E2A0808080010307F7F3010000004067F7F060400;
defparam prom_inst_0.INIT_RAM_07 = 256'h060E1E3E3E1E0E0630383C3E3E3C3830081C3E08083E1C080020202020203C3C;
defparam prom_inst_0.INIT_RAM_08 = 256'h00147F7F147F7F140000070700070700000000065F5F06000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h000000000003070400487A375D4F7A300062660C183066460000123A6B6B2E24;
defparam prom_inst_0.INIT_RAM_0A = 256'h000008083E3E0808082A3E1C1C3E2A080000001C3E63410000000041633E1C00;
defparam prom_inst_0.INIT_RAM_0B = 256'h000103060C183060000000006060000000000808080808080000000060E0A000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000367F494963220000666F49597362000040407F7F424200003E7F4D597F3E;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000070F1971630300003079494B7E3C0000397D4545672700107F7F13161C18;
defparam prom_inst_0.INIT_RAM_0E = 256'h000000006CECA000000000006C6C000000001E3F69494F060000367F49497F36;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000060F595103020000081C3663410000001414141414140000004163361C08;
defparam prom_inst_0.INIT_RAM_10 = 256'h0022634141633E1C00367F49497F7F4100007C7E13137E7C001E1F5D5D417F3E;
defparam prom_inst_0.INIT_RAM_11 = 256'h0072735141633E1C0003011D497F7F410063415D497F7F41001C7F63417F7F41;
defparam prom_inst_0.INIT_RAM_12 = 256'h0063771C087F7F4100013F7F41407030000000417F7F410000007F7F08087F7F;
defparam prom_inst_0.INIT_RAM_13 = 256'h001C3E6341633E1C007F7F180C067F7F007F7F060C067F7F00706040417F7F41;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000327B594D672600466F39197F7F4100005E7F71213F1E00060F09497F7F41;
defparam prom_inst_0.INIT_RAM_15 = 256'h007F7F3018307F7F00001F3F60603F1F00007F7F40407F7F000003417F7F4103;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000041417F7F00007163474D5973670000074F78784F070063771C081C7763;
defparam prom_inst_0.INIT_RAM_17 = 256'h808080808080808000080C0603060C080000007F7F414100006030180C060301;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000286C44447C3800387C44447F3F410040783C545474200000000407030000;
defparam prom_inst_0.INIT_RAM_19 = 256'h00047CF8A4A4BC9800000203497F7E480000185C54547C3800407F3F49487830;
defparam prom_inst_0.INIT_RAM_1A = 256'h00446C38107F7F410000007DFD84C440000000407D7D440000787C04087F7F41;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000387C44447C380000787C04047C7C00787C0C180C7C7C000000407F7F4100;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000247454545C480000181C44787C440084FCF8A4243C1800183C24A4F8FC84;
defparam prom_inst_0.INIT_RAM_1D = 256'h003C7C6030607C3C00001C3C60603C1C00407C3C40407C3C000024447F3E0400;
defparam prom_inst_0.INIT_RAM_1E = 256'h00004141773E08080000644C5C74644C00007CFCA0A0BC9C00446C3810386C44;
defparam prom_inst_0.INIT_RAM_1F = 256'h00787C4643467C780001030203010302000008083E7741410000007777000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h427B7D55557523020000185D57567C3800407A7A40407A3A0000123361E1BF1E;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000143662E2BE1C407A7F55557722000040787C565775200040797D54547521;
defparam prom_inst_0.INIT_RAM_22 = 256'h000001417C7C45010000185C56577D380000195D54547D39021B5D55557D3B02;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000707A2D2D7A700000797D26267D79000000407E7F45000002437D7D450302;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000327B49497B3200497F7F090B7E7C54547C7C5454742000004455577E7C44;
defparam prom_inst_0.INIT_RAM_25 = 256'h004078784243793800407A7B41417B3A000030784A4B79300000327A48487A32;
defparam prom_inst_0.INIT_RAM_26 = 256'h00387C4C54647C3800003D7D40407D3D00397D4444447D3900007AFAA0A0BABA;
defparam prom_inst_0.INIT_RAM_27 = 256'h020B097FFE88C8400000446C38386C44001D3E6749733E5C00206643497F7E68;
defparam prom_inst_0.INIT_RAM_28 = 256'h0040797B424078380000317B4A487830000000417F7E44000040787D57567420;
defparam prom_inst_0.INIT_RAM_29 = 256'h00262F29292F260000282F2F292F260000017B7A33197B7A0001737A0B097B7A;
defparam prom_inst_0.INIT_RAM_2A = 256'h90B9ABEECC1F3F6100003838080808081C22655B4B7D221C00002060454D7830;
defparam prom_inst_0.INIT_RAM_2B = 256'h081C3622081C362222361C0822361C08000060FAFA600000F8D973664C1F3F61;
defparam prom_inst_0.INIT_RAM_2C = 256'h000000FFFF000000FFAAFF55FFAAFF5555AA55AA55AA55AA005500AA005500AA;
defparam prom_inst_0.INIT_RAM_2D = 256'h000070782C2E7B71000072792D2D79720000717B2E2C7870000000FFFF101010;
defparam prom_inst_0.INIT_RAM_2E = 256'h00FCFC04F4F4141400FFFF00FFFF000000FFFF00F7F714141C224155555D221C;
defparam prom_inst_0.INIT_RAM_2F = 256'h000000F0F010101000002B2FFCFC2F2B002424E7E7243C18001F1F1017171414;
defparam prom_inst_0.INIT_RAM_30 = 256'h101010FFFF000000101010F0F01010101010101F1F1010101010101F1F000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0001737A2F2D7B7200417B7E57557722101010FFFF1010101010101010101010;
defparam prom_inst_0.INIT_RAM_32 = 256'h14F4F404F4F41414141717101717141414F4F404FCFC0000141717101F1F0000;
defparam prom_inst_0.INIT_RAM_33 = 256'h00663C3C243C3C6614F7F700F7F71414141414141414141414F7F700FFFF0000;
defparam prom_inst_0.INIT_RAM_34 = 256'h00004555547C7D4500004655557D7D46001C7F63497F7F490000387D57722705;
defparam prom_inst_0.INIT_RAM_35 = 256'h000002457D7D4502000000457F7E44000000000000080E0A00004454567F7D44;
defparam prom_inst_0.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFF101010F0F00000000000001F1F101010000001457C7C4501;
defparam prom_inst_0.INIT_RAM_37 = 256'h0F0F0F0F0F0F0F0F000000447E7F45000000007777000000F0F0F0F0F0F0F0F0;
defparam prom_inst_0.INIT_RAM_38 = 256'h00387C4647457C38003A7D4545457D3A0000143E2A2AFEFC00387C4547467C38;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000081C547E7E42001E3E20207EFE8000397F4647457F3A0001337A4B497B32;
defparam prom_inst_0.INIT_RAM_3A = 256'h00003C7C42437D3C00003A794141793A00003C7D43427C3C00081C14557F7F41;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000103020000000002020202020200000C5D73725C0C000078F9A3A2B8B8;
defparam prom_inst_0.INIT_RAM_3C = 256'hF8D973664C1F35710000282828282828000044445F5F44440000101010101010;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000040C08000000008086B6B0808020359FDA5A5BFDA7F7F017F7F090F06;
defparam prom_inst_0.INIT_RAM_3E = 256'h0010101F1F131200000000101000000000000202000002020000060F090F0600;
defparam prom_inst_0.INIT_RAM_3F = 256'h000000000000000000003C3C3C3C000000001217151D1900000A1F1F15151100;

endmodule //Gowin_pROM
